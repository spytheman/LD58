module main

import gg
import os.asset
import rand
import math

const gwidth = 948
const gheight = 533

enum State {
	working
	paused
	finished
}

@[heap]
struct Game {
mut:
	ctx        &gg.Context = unsafe { nil }
	day        int         = 1
	state      State
	mute_btn   Button
	bins       []Button
	sbin       ?Kind
	day_images []gg.Image
	background gg.Image
	song       &SongPlayer = new_song_player()
	spos       Vec2
	epos       Vec2
	player     Player
	items      []Item
	//
	potential_item_positions []Vec2
}

struct Item {
	pos  Vec2
	img  gg.Image
	kind Kind
}

struct Player {
mut:
	pos    Vec2
	speed  Vec2
	meters u64
	angle  f32
	img    gg.Image
}

fn (mut g Game) restart() {
	g.next_day(g.day)
	g.song.restart()
}

fn (mut g Game) on_mouse(x f32, y f32, e &gg.Event) {
	// eprintln('>> ${@LOCATION}: x: ${x} | y: ${y}')
	g.bins_on_mouse(e)
	if g.mute_btn.clicked(e) {
		g.song.mute()
		g.mute_btn.label = if g.song.mute { 'Unmute' } else { 'Mute' }
	}
}

fn (mut g Game) change_state(nstate State) {
	g.state = nstate
	g.song.pause(nstate == .paused)
}

@[if develop ?]
fn (mut g Game) on_develop(e &gg.Event) {
	if e.typ == .key_down {
		match e.key_code {
			.r { g.restart() }
			.page_up { g.next_day(g.day + 1) }
			.page_down { g.next_day(g.day - 1) }
			else {}
		}
	}
}

fn on_event(e &gg.Event, mut g Game) {
	g.on_develop(e)
	if e.typ == .key_down && e.key_code == .escape {
		g.ctx.quit()
	}
	if e.typ == .char && rune(e.char_code) == `m` {
		g.song.mute()
	}
	if g.state == .finished {
		return
	}
	pause_key := e.key_code in [.space, .p]
	if g.state == .paused && e.typ == .key_up && pause_key {
		g.change_state(.working)
		return
	}
	if g.state == .working && e.typ == .key_up && pause_key {
		g.change_state(.paused)
		return
	}
	if g.state != .working {
		return
	}
	if e.typ == .key_down {
		g.bins_on_key(e)
		match e.key_code {
			.w, .up {
				g.player.speed = Vec2{0, -1}
				g.player.angle = 0
			}
			.s, .down {
				g.player.speed = Vec2{0, 1}
				g.player.angle = math.pi
			}
			.a, .left {
				g.player.speed = Vec2{-1, 0}
				g.player.angle = math.pi / 2
			}
			.d, .right {
				g.player.speed = Vec2{1, 0}
				g.player.angle = -math.pi / 2
			}
			else {}
		}
		return
	}
	x := f32(e.mouse_x)
	y := f32(e.mouse_y)
	g.on_mouse(x, y, e)
}

fn (mut g Game) next_day(nday int) {
	g.day = nday
	if g.day_images.len > 0 {
		lidx := int_max(0, g.day) % g.day_images.len
		g.background = g.day_images[lidx]
	}
	g.find_start_and_exit_spots()
	g.player.speed.zero()
}

fn (mut g Game) player_move() {
	size := 2
	npos := g.player.pos + g.player.speed.mul_scalar(5)
	for y in int(npos.y - size) .. int(npos.y + size) {
		for x in int(npos.x - size) .. int(npos.x + size) {
			c := g.bgpixel(x: x, y: y)
			if c == gg.black {
				return
			}
		}
	}
	g.player.pos = g.player.pos + g.player.speed.mul_scalar(2)
	g.player.meters += u64(g.player.speed.magnitude())
	nc := g.bgpixel(g.player.pos)
	if nc == gg.blue {
		g.next_day(g.day + 1)
	}
	for item_idx, mut item in g.items {
		if g.player.pos.distance(item.pos) < g.player.img.width / 2 {
			g.items.delete(item_idx)
			break
		}
	}
}

fn on_frame(mut g Game) {
	g.song.work() or {}
	g.ctx.begin()
	g.ctx.draw_image(0, 0, g.background.width, g.background.height, g.background)
	for item in g.items {
		g.ctx.draw_rect_filled(item.pos.x, item.pos.y, 5, 5, gg.green)
	}
	g.ctx.draw_image_with_config(
		img_rect: gg.Rect{
			x: g.player.pos.x - g.player.img.width / 2
			y: g.player.pos.y - g.player.img.height / 2
		}
		img:      &g.player.img
		rotation: f32(math.degrees(g.player.angle))
	)
	g.player_move()
	g.bins_draw()
	g.mute_btn.draw(g.ctx)
	g.ctx.draw_text(gwidth - 107, gheight - 34, '${g.state}, day: ${g.day:03}', color: gg.gray)
	g.ctx.draw_text(gwidth - 85, gheight - 18, '${g.player.meters:06}m', color: gg.gray)
	g.ctx.end()
}

fn (mut g Game) bgpixel(pos Vec2) gg.Color {
	x, y := int_max(0, int_min(g.background.width - 1, int(pos.x))), int_max(0, int_min(g.background.height - 1,
		int(pos.y)))
	return unsafe { &gg.Color(g.background.data)[y * g.background.width + x] }
}

fn (mut g Game) find_start_and_exit_spots() {
	g.potential_item_positions.clear()
	g.items.clear()
	g.player.pos.zero()
	g.spos.zero()
	g.epos.zero()
	bp := unsafe { &gg.Color(g.background.data) }
	if isnil(bp) {
		return
	}
	for y in 0 .. gheight {
		for x in 0 .. gwidth {
			c := unsafe { *bp }
			unsafe { bp++ }
			if c.a >= 100 && c.a <= 200 {
				pos := Vec2{x, y}
				_ = pos.str() // TODO: this is needed for tcc, investigate why
				if c.r == 255 {
					g.spos = pos
					g.player.pos = g.spos
				}
				if c.b == 255 {
					g.epos = pos
				}
				if c.g == 255 {
					g.potential_item_positions << pos
				}
			}
		}
	}
	positions := rand.choose(g.potential_item_positions, int_max(5, g.potential_item_positions.len / 5)) or {
		[]
	}
	for ipos in positions {
		g.items << Item{
			pos:  ipos
			kind: unsafe { Kind(rand.int_in_range(0, 4) or { 0 }) }
		}
	}
}

fn main() {
	mut g := &Game{}
	g.mute_btn.pos = Vec2{45, gheight - 16}
	g.mute_btn.size = Vec2{60, 25}
	g.mute_btn.label = 'Mute'
	g.bins_init()
	g.restart()
	g.song.play_ogg_file(asset.get_path('./assets', 'songs/collecting_garbage.ogg'))!
	g.ctx = gg.new_context(
		bg_color:     gg.white
		width:        gwidth
		height:       gheight
		window_title: 'Garbage Collector (LD58)'
		user_data:    g
		frame_fn:     on_frame
		event_fn:     on_event
		font_path:    asset.get_path('./assets', 'fonts/Imprima-Regular.ttf')
		sample_count: 2
	)
	g.player.img = g.ctx.create_image(asset.get_path('./assets', 'images/player.png'))!
	for i in 0 .. 7 + 1 {
		ipath := asset.get_path('./assets', 'images/${i}.png')
		g.day_images << g.ctx.create_image(ipath)!
	}
	g.background = g.day_images[1]
	g.find_start_and_exit_spots()
	g.ctx.run()
}
