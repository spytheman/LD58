module main

#flag wasm32_emscripten -sINITIAL_MEMORY=65536000
#flag wasm32_emscripten --embed-file @DIR/assets/fonts/Imprima-Regular.ttf@/assets/fonts/Imprima-Regular.ttf
#flag wasm32_emscripten --embed-file @DIR/assets/images/0.png@/assets/images/0.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/1.png@/assets/images/1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/2.png@/assets/images/2.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/3.png@/assets/images/3.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/4.png@/assets/images/4.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/5.png@/assets/images/5.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/6.png@/assets/images/6.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/7.png@/assets/images/7.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/glass/cup1.png@/assets/images/items/glass/cup1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/glass/cup2.png@/assets/images/items/glass/cup2.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/glass/cup3.png@/assets/images/items/glass/cup3.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/metal/coin1.png@/assets/images/items/metal/coin1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/metal/coin2.png@/assets/images/items/metal/coin2.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/metal/coin3.png@/assets/images/items/metal/coin3.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/metal/coin4.png@/assets/images/items/metal/coin4.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/organic/apple_bite.png@/assets/images/items/organic/apple_bite.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/organic/leaf1.png@/assets/images/items/organic/leaf1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/organic/remains1.png@/assets/images/items/organic/remains1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/paper/paperball.png@/assets/images/items/paper/paperball.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/paper/sheets1.png@/assets/images/items/paper/sheets1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/paper/toiletroll.png@/assets/images/items/paper/toiletroll.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/plastic/bottle2.png@/assets/images/items/plastic/bottle2.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/plastic/bottle3.png@/assets/images/items/plastic/bottle3.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/plastic/bottle.png@/assets/images/items/plastic/bottle.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/plastic/crap1.png@/assets/images/items/plastic/crap1.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/items/plastic/crap2.png@/assets/images/items/plastic/crap2.png
#flag wasm32_emscripten --embed-file @DIR/assets/images/player.png@/assets/images/player.png
#flag wasm32_emscripten --embed-file @DIR/assets/songs/collecting_garbage.ogg@/assets/songs/collecting_garbage.ogg
